module color_map(
    enemies
);